.title KiCad schematic
.model __Q1 NPN
.model __Q2 NPN
R2 Net-_R1-Pad1_ Net-_Q1-B_ R
R1 Net-_R1-Pad1_ VCC R_Photo
BT1 __BT1
D1 __D1
R3 Net-_Q1-C_ Net-_D2-A_ R
R4 Net-_Q1-C_ Net-_D1-A_ R
Q1 Net-_Q1-C_ Net-_Q1-B_ GND __Q1
M1 __M1
D2 __D2
SW1 __SW1
Q2 VCC Net-_Q2-B_ GND __Q2
R5 Net-_R5-Pad1_ Net-_Q2-B_ R
.end
